shiftreg_inst : shiftreg PORT MAP (
		clock	 => clock_sig,
		shiftin	 => shiftin_sig,
		q	 => q_sig
	);
